// PSW��1 λ״̬�Ĵ���������ֻ�����־λ G��
module psw(
    input  clk,     // ʱ���ź�
    input  g_en,    // ʹ���ź�
    input  g,       // 1 λ����
    output reg gf   // 1 λ���
);

    // ��ʼֵ 0
    initial gf = 1'b0;

    // �� clk �½��أ�g_en = 1 ʱ���� g װ�� gf
    always @(negedge clk) begin
        if (g_en)
            gf <= g;
    end

endmodule