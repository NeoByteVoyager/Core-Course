module controller(
input sm,               // ״̬�ź�
    input [7:0] ir,         // ���ؼ��޸ġ�ֱ������ 8λ IR�������ⲿ���
    input gf,              // ��־λ G
    
  output ld_pc,           
    output in_pc,           
    output [1:0] s,         // RAM��ַѡ��
    output ram_we,          
    output ram_re,          
    output ld_ir,           
    output reg_we,          
    output au_en,           
    output [3:0] ac,        
    output g_en,            
    output in_en,           
    output out_en,          
    output s0,              // �Ĵ���д��Դѡ��
    output sm_en,           
    output [1:0] SR,        
    output [1:0] DR   
);

  
    // 1. ���ָ�� (���ӳ�)
    wire [3:0] opcode = ir[7:4];
    wire [1:0] Rd_raw = ir[3:2];
    wire [1:0] Rs_raw = ir[1:0];

    // 2. ָ������ (���бȽ���)
    localparam MOVA = 4'b0100;
    localparam MOVB = 4'b0101;
    localparam MOVC = 4'b0110;
    localparam MOVD = 4'b0111;
    localparam ADD  = 4'b1000;
    localparam SUB  = 4'b1001;
    localparam JMP  = 4'b1010;
    localparam JG   = 4'b1011;
    localparam IN1  = 4'b1100;
    localparam OUT1 = 4'b1101;
    localparam MOVI = 4'b1110;
    localparam HALT = 4'b1111;

    wire is_mova = (opcode == MOVA);
    wire is_movb = (opcode == MOVB);
    wire is_movc = (opcode == MOVC);
    wire is_movd = (opcode == MOVD);
    wire is_add  = (opcode == ADD);
    wire is_sub  = (opcode == SUB);
    wire is_jmp  = (opcode == JMP);
    wire is_jg   = (opcode == JG);
    wire is_in   = (opcode == IN1);
    wire is_out  = (opcode == OUT1);
    wire is_movi = (opcode == MOVI);
    wire is_halt = (opcode == HALT);

    // 3. ���ٿ����߼�����

    // --- PC ���� ---
    assign ld_pc = sm & (is_jmp | (is_jg & gf));
    assign in_pc = (~sm) | (sm & is_movi);

    // --- RAM ��ַѡ�� (���л��Ż�) ---
    // 00: Fetch/MOVI, 01: MOVC, 10: MOVB
    assign s[0] = sm & is_movc;
    assign s[1] = sm & is_movb;

    // --- RAM ��д ---
    assign ram_re = (~sm) | (sm & (is_movc | is_movi));
    assign ram_we = sm & is_movb;

    // --- �Ĵ������� ---
    assign s0 = ~(sm & is_movd); // ֻ�� MOVD ʱΪ 0������Ϊ 1

    assign reg_we = sm & (is_mova | is_movc | is_movd | is_add | is_sub | is_in | is_movi);

    // Ѱַ�߼��Ż�
    assign SR = (is_jmp | is_jg | is_movd) ? 2'b11 : Rs_raw;
    
    // �����Ƕ�� MUX �ۺ���ͨ������úܺ�
    assign DR = is_movi ? 2'b00 : (is_movd ? 2'b11 : Rd_raw);

    // --- AU ���� ---
    assign au_en = sm & (is_mova | is_add | is_sub | is_out | is_movb);
    
    // ac �����߼�ֱ�ۼ���
    assign ac = (is_add) ? 4'b1000 : 
                (is_sub) ? 4'b1001 : 
                (is_mova | is_out | is_movb) ? 4'b0100 : 4'b0000;

    // --- ���� ---
    assign sm_en  = ~(sm & is_halt);
    assign ld_ir  = ~sm;
    assign g_en   = sm & is_sub;
    assign in_en  = sm & is_in;
    assign out_en = sm & is_out;

endmodule