module reg_group (
    input wire clk,
    input wire we,
    input wire [1:0] sr,
    input wire [1:0] dr,
    input wire [7:0] i,
    output reg [7:0] s,
    output reg [7:0] d
);

    // 4��8λ�Ĵ���
    reg [7:0] R0, R1, R2, R3;
    initial begin
        R0 = 8'h01;
        R1 = 8'b0000_0000;
        R2 = 8'b0000_0000;
        R3 = 8'h07;
    end
    
      // ������������߼���S�ڣ�
	always @(*) begin
		case (sr)
			2'b00: s = R0;
			2'b01: s = R1;
			2'b10: s = R2;
			2'b11: s = R3;
			default: s = 8'b0; // ��ֹ����
		endcase
	end

	// ������������߼���D�ڣ�
	always @(*) begin
		case (dr)
			2'b00: d = R0;
			2'b01: d = R1;
			2'b10: d = R2;
			2'b11: d = R3;
			default: d = 8'b0;
		endcase
	end
    
    // д������ʱ���½��ش���
    always @(negedge clk) begin
        if (we) begin
            case (dr)
                2'b00: R0 <= i;
                2'b01: R1 <= i;
                2'b10: R2 <= i;
                2'b11: R3 <= i;
            endcase
        end
    end
    
	 


endmodule