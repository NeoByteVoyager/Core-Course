module half_adder(
S,I,Y	
);
input [1:0]S;
input [3:0]I;
output Y;
reg Y;
always @(S or Y)
begin
case(S)
2'b00:Y=I[0];
2'b01:Y=I[1];
2'b10:Y=I[2];
2'b11:Y=I[3];
default:Y=1'bx;
endcase
end
endmodule 