module sm (
    input wire clk,
    input wire sm_en,
    output reg [1:0] sm // ���޸ġ������Ϊ 2 λ��
);
    // ����״̬���ƣ������Ķ�
    parameter S_FETCH = 2'b00;
    parameter S_PREP  = 2'b01;
    parameter S_EXEC  = 2'b10;

    initial sm = S_FETCH;
    
    // �����½��ش��������Buffer������������
    always @(negedge clk) begin
        if (sm_en) begin
            case (sm)
                S_FETCH: sm <= S_PREP;
                S_PREP:  sm <= S_EXEC;
                S_EXEC:  sm <= S_FETCH;
                default: sm <= S_FETCH;
            endcase
        end
    end
endmodule