// IR��8 λָ��Ĵ���
module ir(
    input        clk,    // ʱ���ź�
    input        ld_ir,  // װ��ʹ���ź�
    input  [7:0] a,      // 8 λ����
    output reg [7:0] x   // 8 λ���
);

    // ��ʼֵ 00000000
    initial x = 8'b00000000;

    // �� clk �½��أ�ld_ir = 1 ʱ�������� a װ��Ĵ���
    always @(negedge clk) begin
        if (ld_ir)
            x <= a;
    end

endmodule