module controller(
    input sm,               // ״̬�źţ�0Ϊȡָ��1Ϊִ��
    input mova, movb, movc, movd, add, sub, jmp, jg, in1, out1, movi, halt, // ���������
    input gf,               // ״̬�Ĵ�����־λ G
    output ld_pc,           // ����PC
    output in_pc,           // PC����
    output s1, s2,          // RAM��ַѡ��
    output ram_we,          // RAMдʹ�� (WR)
    output ram_re,          // RAM��ʹ�� (RE)
    output ld_ir,           // ָ��Ĵ���װ��
    output reg_we,          // ͨ�üĴ�����дʹ��
    output au_en,           // ���㵥Ԫ���ʹ��
    output [3:0] ac,        // ���㵥Ԫ���ܿ���
    output g_en,            // ״̬�Ĵ���дʹ��
    output in_en,           // �����豸ʹ��
    output out_en,          // ����豸ʹ��
    output s0,              // �Ĵ�������������Դѡ�� (0:PC, 1:����)
    output sm_en            // ״̬����תʹ��
);

    // 1. PC �����߼�
    // ��ת�߼���ִ�н׶�(sm=1) �� (��������ת �� ��������ת��G=1)
    assign ld_pc = sm & (jmp | (jg & gf));
    // �����߼���ȡָ�׶�(sm=0)
    assign in_pc = ~sm;

    // 2. RAM ��ַѡ���߼� (s2, s1)
    // 00: PC(ȡָ), 01: S��(movc), 10: D��(movb)
    assign s1 = sm & movc;
    assign s2 = sm & movb;

    // 3. RAM ��д�߼�
    assign ram_we = sm & movb;         // ִ��movbʱд��RAM
    assign ram_re = (~sm) | (sm & movc); // ȡָ�� �� ִ��movcʱ��ȡ

    // 4. IR װ���߼�
    assign ld_ir = ~sm;                // ����ȡָ��װ��

    // 5. ͨ�üĴ�����д���߼� (reg_we)
    // �����޸�Ŀ�ļĴ�����ָ���Ҫдʹ��
    assign reg_we = sm & (mova | movc | movd | add | sub | in1 | movi);

    // 6. ���㵥Ԫ���� (AU)
    // AU��Ҫ��������ߵ�ָ��
    assign au_en = sm & (mova | add | sub | out1);
    // AU������ӳ��
    assign ac = add ? 4'b1000 : 
               (sub ? 4'b1001 : 
               (mova ? 4'b0100 : 4'b0000));

    // 7. ״̬λ���� (G_EN)
    assign g_en = sm & sub;            // ������ָ�����G��־

    // 8. ����/����豸ʹ��
    assign in_en = sm & in1;
    assign out_en = sm & out1;

    // 9. �Ĵ�����������Դѡ�� (s0)
    // 0: ����PC (movd), 1: �������� (����ָ��)
    assign s0 = ~(sm & movd);

    // 10. ͣ������
    assign sm_en = ~halt;              // halt��Чʱ��ֹSM��ת��ϵͳֹͣ

endmodule