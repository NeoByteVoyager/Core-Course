module pc(
    input        clk,    // ʱ��
    input        ld_pc,  // װ�ؿ���
    input        in_pc,  // ��������
    input  [7:0] a,      // 8 λ���루��ת��ַ��
    output reg [7:0] c   // 8 λ�������ǰ PC��
);

    initial c = 8'b00000000;   // ��ʼȡֵΪ 0����һ��ָ���ַ��

    always @(negedge clk) begin
        if (ld_pc)
            c <= a;              // װ����ת��ַ
        else if (in_pc)
            c <= c + 8'b00000001; // ˳��ִ�У��Լ� 1
        // ���򱣳ֲ���
    end

endmodule