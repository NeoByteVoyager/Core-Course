module controller(
    input [1:0] sm,         // ״̬�źű�Ϊ2λ��00ȡָ��01׼����10ִ��
    input mova, movb, movc, movd, add, sub, jmp, jg, in1, out1, movi, halt, 
    input [7:0] ir,     
    input gf,               

    output ld_pc, in_pc,
    output  [1:0]s,
    output ram_re, ram_we, ld_dr, ld_ir, reg_we, s0,
    output [1:0]  SR, DR,
    
    output  au_en, 
    output [3:0] ac,
    output g_en,in_en, out_en, sm_en,
    output decoder_en
    
);
	
	

    wire fetch = (sm == 2'b00);
    wire prep  = (sm == 2'b01);
    wire exec  = (sm == 2'b10);
    
   
   
	assign in_pc  = fetch | (exec & movi);
    assign ld_pc  = exec & (jmp | (jg & gf));
    
   
    assign s = exec  ? (movc ? 2'b01 :  
                        movb ? 2'b10 :  
                        2'b00) :        
               2'b00;


    assign ram_re = fetch | (exec & (movc | movi)); 
    assign ram_we = exec & movb;
	
	assign ld_ir  = fetch;
	
	assign decoder_en = sm[0] | sm[1];//
	
    assign ld_dr  = prep; // DR ��Ȼ��׼�����ڹ���������Ƕ����ڵ�֤��
    
	assign s0     = (exec & movd) ? 1'b0 : 1'b1;//
    assign reg_we = exec & (mova | movc | movd | add | sub | in1 | movi);
    
    assign SR     = ir[1:0];
    assign DR     = ir[3:2];
    
    assign au_en  = exec & (mova | add | sub | movb | out1);//
    assign ac     = ir[7:4];
    assign g_en   = exec & sub;
    
    assign in_en  = exec & in1;
    assign out_en = exec & out1;
    
    
	assign sm_en  = ~(exec & halt);
endmodule